module rename(
	input  logic       clk,
	input  logic       rst_ni,
	input  br_result_t br_result_i,
	input  p_reg_t     p_commit_i,   //in-order commit
	input  dinstr_t    dinstr_i,
	output rinstr_t    rinstr_o,
	output logic       rn_full_o
);

	/* Your Code Here */
	//...
	//...
	//...

endmodule
